
// 8 bit number //

interface number;
    logic [7:0] bits;
endinterface

// 4 bit address //

interface address;
    logic [3:0] bits;
endinterface

